module write_back (/* create ports Here */);

endmodule
