module memory (/* Create Ports Here */);


endmodule
