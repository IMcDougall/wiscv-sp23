module fetch ( /*Create Ports Here */);



endmodule
