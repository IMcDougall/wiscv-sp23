module execute (/* create Ports Here*/);

endmodule
