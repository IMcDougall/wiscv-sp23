module decode (/* create Ports Here*/);


endmodule
