module register_file (/* Create Ports Here*/);



endmodule
